** Generated for: hspiceD
** Generated on: Oct 26 11:33:46 2022
** Design library name: ELEC402
** Design cell name: buffer
** Design view name: schematic
.GLOBAL vdd!


.PROBE TRAN
+    V(in)
+    V(out)
.TRAN 200e-15 2e-9 START=0.0

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.LIB "/ubc/ece/data/cmc2/kits/ncsu_pdk/FreePDK15/hspice/models/fet.inc" CMG

** Library name: ELEC402
** Cell name: buffer
** View name: schematic
m0 vdd! in out vdd! nfet AD=608e-18 AS=608e-18 PD=168e-9 PS=168e-9 M=2
m1 0 in out 0 pfet AD=608e-18 AS=608e-18 PD=168e-9 PS=168e-9 M=2
c0 out 0 1e-15
v0 in 0 PWL 0 0 500e-12 0 1e-9 900e-3 1.5e-9 0 TD=0
.END
